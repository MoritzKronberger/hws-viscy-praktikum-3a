----------------------------------------------------------------------------------------
-- This file is part of the VISCY project.
-- (C) 2007-2021 Gundolf Kiefer, Fachhochschule Augsburg, University of Applied Sciences
-- (C) 2018 Michael Schäferling, Hochschule Augsburg, University of Applied Sciences
--
-- Description:
-- This is a testbench for the VISCY CPU
----------------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity CPU_TB is
end CPU_TB;


architecture TESTBENCH of CPU_TB is
    -- Declare CPU component (Unit Under Test - UUT)
    component CPU is
        port (
            clk:    in    std_logic;                      -- clock signal
            reset:  in    std_logic;                      -- reset CPU
            adr:    out   std_logic_vector (15 downto 0); -- memory address
            rdata:  in    std_logic_vector (15 downto 0); -- data read from memory
            wdata:  out   std_logic_vector (15 downto 0); -- data to write to memory
            rd:     out   std_logic;                      -- read from memory
            wr:     out   std_logic;                      -- write to memory
            ready:  in    std_logic                       -- ready signal
            );
        end component;

    -- Point CPU component to the submodule's RTL architecture
    for UUT: CPU use entity WORK.CPU(RTL);

    -- Internal signals
    signal clk:   std_logic := '0';              -- clock signal
    signal reset: std_logic := '0';              -- reset CPU
    signal ready: std_logic := '0';              -- ready signal
    signal adr:   std_logic_vector(15 downto 0); -- memory address
    signal rdata: std_logic_vector(15 downto 0); -- data read from memory
    signal wdata: std_logic_vector(15 downto 0); -- data to write to memory
    signal rd:    std_logic;                     -- read from memory
    signal wr:    std_logic;                     -- write to memory

    -- Internal constants
    constant clk_period: time := 10 ns;
    constant mem_delay: time := 25 ns;

    -- Memory content (generated by viscy2l)
    type t_memory is array (0 to 42) of std_logic_vector (15 downto 0);
    signal mem_content: t_memory := (
        16#0000# => "0011000000000000",  --        xor r0, r0, r0 ; r0 := 00000000 00000000 (=0) | Funktioniert nicht, da Bits = 'U'?
        16#0001# => "0011011111111100",  --        xor r7, r7, r7 ; r7 := 00000000 00000000 (=0) | Funktioniert nicht, da Bits = 'U'?
        16#0002# => "0100000100000101",  --        ldil r1, 5     ; r1 := 00000000 00000101 (lo=5)
        16#0003# => "0100101000001000",  --        ldih r2, 8       ; r2 := 00001000 00000000 (2048)
        16#0004# => "0100001100000110",  --        ldil r3, 6       ; r3 := -------- 00000110 (lo=6)
        16#0005# => "0100101100001100",  --        ldih r3, 12      ; r3 := 00001100 00000110 (=3078)
        16#0006# => "0100000100001010",  --        ldil r1, 10 ; r1 := -------- 00001010 (lo=10)
        16#0007# => "0100100100000000",  --        ldih r1, 0  ; r1 := 00000000 00001010 (=10)
        16#0008# => "0100001000000010",  --        ldil r2, 2  ; r2 := -------- 00000010 (lo=2)
        16#0009# => "0100101000010001",  --        ldih r2, 17 ; r2 := 00010001 00000010 (=4354)
        16#000a# => "0000010000101000",  --        add r4, r1, r2   ; r4 := 00010001 00001100 (=4364)
        16#000b# => "0100011100001100",  --        ldil r7, 0x0C
        16#000c# => "0100111100010001",  --        ldih r7, 0x11  ; r7 := 00010001 00001100 (=4364)
        16#000d# => "0011000010011100",  --        xor r0, r4, r7 ; r0 := 00000000 00000000 (0)
        16#000e# => "0000110101000100",  --        sub r5, r2, r1   ; r5 := 00010000 11111000 (=4344)
        16#000f# => "0100011111111000",  --        ldil r7, 0xF8
        16#0010# => "0100111100010000",  --        ldih r7, 0x10  ; r7 := 00010000 11111000 (=4344)
        16#0011# => "0011000010111100",  --        xor r0, r5, r7 ; 00000000 00000000 (0)
        16#0012# => "0001011001000000",  --        sal r6, r2       ; r6 := 00100010 00000100 (=8708)
        16#0013# => "0100011100000100",  --        ldil r7, 0x04
        16#0014# => "0100111100100010",  --        ldih r7, 0x22  ; r7 := 00100010 00000100 (=8708)
        16#0015# => "0011000011011100",  --        xor r0, r6, r7 ; r0 := 00000000 00000000 (0)
        16#0016# => "0001101101000000",  --        sar r3, r2       ; r3 := 00001000 10000001 (=2177)
        16#0017# => "0100011110000001",  --        ldil r7, 0x81
        16#0018# => "0100111100001000",  --        ldih r7, 0x08  ; r7 := 00001000 10000001 (=2177)
        16#0019# => "0011000001111100",  --        xor r0, r3, r7 ; r0 := 00000000 00000000 (0)
        16#001a# => "0010001100101000",  --        and r3, r1, r2 ; r3 := 00000000 00000010 (=2)
        16#001b# => "0100011100000010",  --        ldil r7, 0x02
        16#001c# => "0100111100000000",  --        ldih r7, 0x00  ; r7 := 00000000 00000010 (=2)
        16#001d# => "0011000001111100",  --        xor r0, r3, r7 ; r0 := 00000000 00000000 (0)
        16#001e# => "0010101100101000",  --        or r3, r1, r2    ; r3 := 00010001 00001010 (=4362)
        16#001f# => "0100011100001010",  --        ldil r7, 0x0A
        16#0020# => "0100111100010001",  --        ldih r7, 0x11  ; r7 := 00010001 00001010 (=4362)
        16#0021# => "0011000001111100",  --        xor r0, r3, r7 ; r0 := 00000000 00000000 (0)
        16#0022# => "0011001100101000",  --        xor r3, r1, r2   ; r3 := 00010001 00001000 (=4360)
        16#0023# => "0100011100001000",  --        ldil r7, 0x08
        16#0024# => "0100111100010001",  --        ldih r7, 0x11  ; r7 := 00010001 00001000 (=4360)
        16#0025# => "0011000001111100",  --        xor r0, r3, r7 ; r0 := 00000000 00000000 (0)
        16#0026# => "0011101101000000",  --        not r3, r2        ; r3 := 11101110 11111101 (=61181)
        16#0027# => "0100011111111101",  --        ldil r7, 0xFD
        16#0028# => "0100111111101110",  --        ldih r7, 0xEE  ; r7 := 11101110 11111101 (=61181)
        16#0029# => "0011000001111100",  --        xor r0, r3, r7 ; 00000000 00000000 (0)
        16#002a# => "1000100000000000",  --        halt ; Prozessor anhalten
        others => "UUUUUUUUUUUUUUUU"
    );

BEGIN
    -- Instantiate the CPU (UUT)
    UUT: CPU port map (
            clk => clk,
            reset => reset,
            adr => adr,
            rdata => rdata,
            wdata => wdata,
            rd => rd,
            wr => wr,
            ready => ready
         );

    -- Process to simulate the memory behavior
    memory: process
    begin
        -- Disable ready
        ready <= '0';
        -- Wait until CPU wants to read or write
        wait on rd, wr;
        -- In read mode
        if rd = '1' then
            wait for mem_delay; -- simulate memory delay
            -- Set read-data from memory-address-data
            if is_x (adr) then
                rdata <= (others => 'X'); -- fill read-data with X if memory address is X
            else
                rdata <= mem_content (to_integer (unsigned (adr))); -- otherwise, load memory content from memory address into read-data
            end if;
            -- Enable ready (data can now be used by CPU)
            ready <= '1';
            -- Wait until CPU disables read mode
            wait until rd = '0';
            -- Fill read-data with X (invalid data, which should not be used by CPU since rd = 0)
            rdata <= (others => 'X');
            wait for mem_delay; -- simulate memory delay
            -- Disable ready
            ready <= '0';
        -- In write mode
        elsif wr = '1' then
            wait for mem_delay; -- simulate memory delay
            -- Set memory-address-data from write-data (if address is not X)
            if not is_x(adr) then
                mem_content (to_integer (unsigned (adr))) <= wdata;
            end if;
            -- Enable ready (write was successful)
            ready <= '1';
            -- Wait until CPU disables write mode
            wait until wr = '0';
            wait for mem_delay; -- simulate memory delay
            -- Disable ready
            ready <= '0';
        end if;
    end process;


  -- Main testbench process
  testbench: process
    
    procedure run_cycle is
    begin
      clk <= '0';
      wait for clk_period / 2;
      clk <= '1';
      wait for clk_period / 2;
    end procedure;

    -- End testbench after n cycles without read signal
    variable read_tb_timeout: integer := 20;
    
  begin

    -- Reset CPU on startup
    reset <= '1';
    run_cycle;
    reset <= '0';

    -- Run clock cycles
    -- Exit loop if read timeout expires
    L: while read_tb_timeout > 0 loop
        run_cycle;
        -- Increment timeout if read signal is not set
        IF rd = '0' THEN
            read_tb_timeout := read_tb_timeout - 1;
        END IF;
    end loop;
    
    -- Print a note & finish simulation now
    assert false report "Simulation finished" severity note;
    wait; -- wait forever (stop simulation)

  end process;

end architecture;
