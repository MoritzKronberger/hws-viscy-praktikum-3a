----------------------------------------------------------------------------------------
-- This file is part of the VISCY project.
-- (C) 2007-2021 Gundolf Kiefer, Fachhochschule Augsburg, University of Applied Sciences
-- (C) 2018 Michael Schäferling, Hochschule Augsburg, University of Applied Sciences
--
-- Description:
-- This is a testbench for the VISCY CPU
----------------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity CPU_TB is
end CPU_TB;


architecture TESTBENCH of CPU_TB is
    -- Declare CPU component (Unit Under Test - UUT)
    component CPU is
        port (
            clk:    in    std_logic;                      -- clock signal
            reset:  in    std_logic;                      -- reset CPU
            adr:    out   std_logic_vector (15 downto 0); -- memory address
            rdata:  in    std_logic_vector (15 downto 0); -- data read from memory
            wdata:  out   std_logic_vector (15 downto 0); -- data to write to memory
            rd:     out   std_logic;                      -- read from memory
            wr:     out   std_logic;                      -- write to memory
            ready:  in    std_logic                       -- ready signal
            );
        end component;

    -- Point CPU component to the submodule's RTL architecture
    for UUT: CPU use entity WORK.CPU(RTL);

    -- Internal signals
    signal clk:   std_logic := '0';              -- clock signal
    signal reset: std_logic := '0';              -- reset CPU
    signal ready: std_logic := '0';              -- ready signal
    signal adr:   std_logic_vector(15 downto 0); -- memory address
    signal rdata: std_logic_vector(15 downto 0); -- data read from memory
    signal wdata: std_logic_vector(15 downto 0); -- data to write to memory
    signal rd:    std_logic;                     -- read from memory
    signal wr:    std_logic;                     -- write to memory

    -- Internal constants
    constant clk_period: time := 10 ns;
    constant mem_delay: time := 25 ns;

    -- Memory content (generated by viscy2l) ...
    type t_memory is array (0 to 272) of std_logic_vector (15 downto 0);
    signal mem_content: t_memory := (
        16#0000# => "0100000000000000",  --         ldil r0, result & 255
        16#0001# => "0100100000000001",  --         ldih r0, result >> 8 ; r0 := result (Adresse)
        16#0002# => "0100000100000001",  --         ldil r1, 1           ; r1 := --------00000001 (lo=1)
        16#0003# => "0100100100000000",  --         ldih r1, 0           ; r1 := 0000000000000001 (=1)
        16#0004# => "0100001000000101",  --         ldil r2, 5     ; r0 = --------00000101 (lo=5)
        16#0005# => "0101100000001000",  --         st [r0], r2    ; Ergebnis schreiben
        16#0006# => "0000000000000100",  --         add r0, r0, r1 ; Zieladresse inkrementieren
        16#0007# => "0100101100001000",  --         ldih r3, 8     ; r3 = 00001000-------- (hi=8)
        16#0008# => "0101100000001100",  --         st [r0], r3    ; Ergebnis schreiben
        16#0009# => "0000000000000100",  --         add r0, r0, r1 ; Zieladresse inkrementieren
        16#000a# => "0100010000000110",  --         ldil r4, 6     ; r4 := --------00000110 (lo=6)
        16#000b# => "0100110000001100",  --         ldih r4, 12    ; r4 := 0000110000000110 (=3078)
        16#000c# => "0101100000010000",  --         st [r0], r4    ; Ergebnis schreiben
        16#000d# => "0000000000000100",  --         add r0, r0, r1 ; Zieladresse inkrementieren
        16#000e# => "0000110100000100",  --         sub r5, r0, r1 ; letzte Zieladresse erhalten
        16#000f# => "0101011010100000",  --         ld r6, [r5]
        16#0010# => "0101100000011000",  --         st [r0], r6    ; Ergebnis schreiben
        16#0011# => "0000000000000100",  --         add r0, r0, r1 ; Zieladresse inkrementieren
        16#0012# => "0100010100001010",  --         ldil r5, 10 ; r5 := --------00001010 (lo=10)
        16#0013# => "0100110100000000",  --         ldih r5, 0  ; r5 := 0000000000001010 (=10)
        16#0014# => "0100011000000010",  --         ldil r6, 2  ; r6 := --------00000010 (lo=2)
        16#0015# => "0100111000010001",  --         ldih r6, 17 ; r6 := 0001000100000010 (=4354)
        16#0016# => "0011011111111100",  --         xor r7, r7, r7 ; r7 := 0000000000000000 (=0)
        16#0017# => "0000011110111000",  --         add r7, r5, r6 ; r7 := 0001000100001100 (=4364)
        16#0018# => "0101100000011100",  --         st [r0], r7    ; Ergebnis schreiben
        16#0019# => "0000000000000100",  --         add r0, r0, r1 ; Zieladresse inkrementieren
        16#001a# => "0011011111111100",  --         xor r7, r7, r7 ; r7 := 0000000000000000 (=0)
        16#001b# => "0000111111010100",  --         sub r7, r6, r5 ; r7 := 0001000011111000 (=4344)
        16#001c# => "0101100000011100",  --         st [r0], r7    ; Ergebnis schreiben
        16#001d# => "0000000000000100",  --         add r0, r0, r1 ; Zieladresse inkrementieren
        16#001e# => "0011011111111100",  --         xor r7, r7, r7 ; r7 := 0000000000000000 (=0)
        16#001f# => "0001011111000000",  --         sal r7, r6     ; r7 := 0010001000000100 (=8708)
        16#0020# => "0101100000011100",  --         st [r0], r7    ; Ergebnis schreiben
        16#0021# => "0000000000000100",  --         add r0, r0, r1 ; Zieladresse inkrementieren
        16#0022# => "0011011111111100",  --         xor r7, r7, r7 ; r7 := 0000000000000000 (=0)
        16#0023# => "0001111111000000",  --         sar r7, r6     ; r7 := 0000100010000001 (=2177)
        16#0024# => "0101100000011100",  --         st [r0], r7    ; Ergebnis schreiben
        16#0025# => "0000000000000100",  --         add r0, r0, r1 ; Zieladresse inkrementieren
        16#0026# => "0011011111111100",  --         xor r7, r7, r7 ; r7 := 0000000000000000 (=0)
        16#0027# => "0010011110111000",  --         and r7, r5, r6 ; r7 := 0000000000000010 (=2)
        16#0028# => "0101100000011100",  --         st [r0], r7    ; Ergebnis schreiben
        16#0029# => "0000000000000100",  --         add r0, r0, r1 ; Zieladresse inkrementieren
        16#002a# => "0011011111111100",  --         xor r7, r7, r7 ; r7 := 0000000000000000 (=0)
        16#002b# => "0010111110111000",  --         or r7, r5, r6  ; r7 := 0001000100001010 (=4362)
        16#002c# => "0101100000011100",  --         st [r0], r7    ; Ergebnis schreiben
        16#002d# => "0000000000000100",  --         add r0, r0, r1 ; Zieladresse inkrementieren
        16#002e# => "0011011111111100",  --         xor r7, r7, r7 ; r7 := 0000000000000000 (=0)
        16#002f# => "0011011110111000",  --         xor r7, r5, r6 ; r7 := 0001000100001000 (=4360)
        16#0030# => "0101100000011100",  --         st [r0], r7    ; Ergebnis schreiben
        16#0031# => "0000000000000100",  --         add r0, r0, r1 ; Zieladresse inkrementieren
        16#0032# => "0011011111111100",  --         xor r7, r7, r7 ; r7 := 0000000000000000 (=0)
        16#0033# => "0011111111000000",  --         not r7, r6     ; r7 := 1110111011111101 (=61181)
        16#0034# => "0101100000011100",  --         st [r0], r7    ; Ergebnis schreiben
        16#0035# => "0000000000000100",  --         add r0, r0, r1 ; Zieladresse inkrementieren
        16#0036# => "0100001000000100",  --         ldil r2, 4              ; r2 := --------00000100 (lo=4)
        16#0037# => "0100101000000000",  --         ldih r2, 0              ; r2 := 0000000000000100 (=4)
        16#0038# => "0100001100111101",  --         ldil r3, jumpskip & 255
        16#0039# => "0100101100000000",  --         ldih r3, jumpskip >> 8 ; r3 := jumpskip (Adresse)
        16#003a# => "1000000001100000",  --         jmp r3                 ; jump to jumpskip label
        16#003b# => "0100001011111111",  --         ldil r2, 0xFF          ; should be skipped
        16#003c# => "0100101011111111",  --         ldih r2, 0xFF          ; should be skipped
        16#003d# => "0101100000001000",  --         st [r0], r2            ; Ergebnis schreiben
        16#003e# => "0000000000000100",  --         add r0, r0, r1         ; Zieladresse inkrementieren
        16#003f# => "0100001000001011",  --         ldil r2, 11            ; r2 := --------00001011 (lo=11)
        16#0040# => "0100101000110100",  --         ldih r2, 52            ; r2 := 0011010000001011 (=13323)
        16#0041# => "0011010010010000",  --         xor r4, r4, r4
        16#0042# => "0100001101000111",  --         ldil r3, jztskip & 255
        16#0043# => "0100101100000000",  --         ldih r3, jztskip >> 8 ; r3 := jztskip (Adresse)
        16#0044# => "1001000001110000",  --         jz r4, r3             ; jump to jztskip label
        16#0045# => "0100001011111111",  --         ldil r2, 0xFF         ; should be skipped
        16#0046# => "0100101011111111",  --         ldih r2, 0xFF         ; should be skipped
        16#0047# => "0101100000001000",  --         st [r0], r2           ; Ergebnis schreiben
        16#0048# => "0000000000000100",  --         add r0, r0, r1        ; Zieladresse inkrementieren
        16#0049# => "0100001011111111",  --         ldil r2, 0xFF         ; r2 := --------11111111
        16#004a# => "0100101011111111",  --         ldih r2, 0xFF         ; r2 := 1111111111111111
        16#004b# => "0100010000000001",  --         ldil r4, 1            ; r4 := --------00000001 (lo=1)
        16#004c# => "0100001101010001",  --         ldil r3, jzfskip & 255
        16#004d# => "0100101100000000",  --         ldih r3, jzfskip >> 8 ; r3 := jzfskip (Adresse)
        16#004e# => "1001000001110000",  --         jz r4, r3             ; do not jump to jzfskip label
        16#004f# => "0100001000010001",  --         ldil r2, 17           ; should be executed, r2 := --------00010001 (lo=17)
        16#0050# => "0100101000010111",  --         ldih r2, 23           ; should be executed, r2 := 0001011100010001 (=5905)
        16#0051# => "0101100000001000",  --         st [r0], r2           ; Ergebnis schreiben
        16#0052# => "0000000000000100",  --         add r0, r0, r1        ; Zieladresse inkrementieren
        16#0053# => "0100001000101111",  --         ldil r2, 47            ; r2 := --------00101111 (lo=47)
        16#0054# => "0100101000110100",  --         ldih r2, 52            ; r2 := 0011010000101111 (=13359)
        16#0055# => "0100010000000001",  --         ldil r4, 1             ; r4 := --------00000001 (lo=1)
        16#0056# => "0100001101011011",  --         ldil r3, jnztskip & 255
        16#0057# => "0100101100000000",  --         ldih r3, jnztskip >> 8 ; r3 := jnztskip (Adresse)
        16#0058# => "1001100001110000",  --         jnz r4, r3             ; jump to jnztskip label
        16#0059# => "0100001011111111",  --         ldil r2, 0xFF          ; should be skipped
        16#005a# => "0100101011111111",  --         ldih r2, 0xFF          ; should be skipped
        16#005b# => "0101100000001000",  --         st [r0], r2            ; Ergebnis schreiben
        16#005c# => "0000000000000100",  --         add r0, r0, r1         ; Zieladresse inkrementieren
        16#005d# => "0100001011111111",  --         ldil r2, 0xFF          ; r2 := --------11111111
        16#005e# => "0100101011111111",  --         ldih r2, 0xFF          ; r2 := 1111111111111111
        16#005f# => "0011010010010000",  --         xor r4, r4, r4         ; r4 := 0000000000000000 (=0)
        16#0060# => "0100001101100101",  --         ldil r3, jnzfskip & 255
        16#0061# => "0100101100000000",  --         ldih r3, jnzfskip >> 8 ; r3 := jnzfskip (Adresse)
        16#0062# => "1001100001110000",  --         jnz r4, r3             ; do not jump to jnzfskip label
        16#0063# => "0100001000001000",  --         ldil r2, 8             ; should be executed, r2 := --------00001000 (lo=8)
        16#0064# => "0100101000010000",  --         ldih r2, 16            ; should be executed, r2 := 0001000000001000 (=4104)
        16#0065# => "0101100000001000",  --         st [r0], r2            ; Ergebnis schreiben
        16#0066# => "0000000000000100",  --         add r0, r0, r1         ; Zieladresse inkrementieren
        16#0067# => "1000100000000000",  --         halt ; Prozessor anhalten
        16#0100# => "0000000000000000",  -- result: .res 17 ; 17 Worte reservieren (für alle Test-Cases)
        16#0101# => "0000000000000000",
        16#0102# => "0000000000000000",
        16#0103# => "0000000000000000",
        16#0104# => "0000000000000000",
        16#0105# => "0000000000000000",
        16#0106# => "0000000000000000",
        16#0107# => "0000000000000000",
        16#0108# => "0000000000000000",
        16#0109# => "0000000000000000",
        16#010a# => "0000000000000000",
        16#010b# => "0000000000000000",
        16#010c# => "0000000000000000",
        16#010d# => "0000000000000000",
        16#010e# => "0000000000000000",
        16#010f# => "0000000000000000",
        16#0110# => "0000000000000000",
        others => "UUUUUUUUUUUUUUUU"
    );

BEGIN
    -- Instantiate the CPU (UUT)
    UUT: CPU port map (
            clk => clk,
            reset => reset,
            adr => adr,
            rdata => rdata,
            wdata => wdata,
            rd => rd,
            wr => wr,
            ready => ready
         );

    -- Process to simulate the memory behavior
    memory: process
    begin
        -- Disable ready
        ready <= '0';
        -- Wait until CPU wants to read or write
        wait on rd, wr;
        -- In read mode
        if rd = '1' then
            wait for mem_delay; -- simulate memory delay
            -- Set read-data from memory-address-data
            if is_x (adr) then
                rdata <= (others => 'X'); -- fill read-data with X if memory address is X
            else
                rdata <= mem_content (to_integer (unsigned (adr))); -- otherwise, load memory content from memory address into read-data
            end if;
            -- Enable ready (data can now be used by CPU)
            ready <= '1';
            -- Wait until CPU disables read mode
            wait until rd = '0';
            -- Fill read-data with X (invalid data, which should not be used by CPU since rd = 0)
            rdata <= (others => 'X');
            wait for mem_delay; -- simulate memory delay
            -- Disable ready
            ready <= '0';
        -- In write mode
        elsif wr = '1' then
            wait for mem_delay; -- simulate memory delay
            -- Set memory-address-data from write-data (if address is not X)
            if not is_x(adr) then
                mem_content (to_integer (unsigned (adr))) <= wdata;
            end if;
            -- Enable ready (write was successful)
            ready <= '1';
            -- Wait until CPU disables write mode
            wait until wr = '0';
            wait for mem_delay; -- simulate memory delay
            -- Disable ready
            ready <= '0';
        end if;
    end process;


  -- Main testbench process
  testbench: process
    
    procedure run_cycle is
    begin
      clk <= '0';
      wait for clk_period / 2;
      clk <= '1';
      wait for clk_period / 2;
    end procedure;

    -- End testbench after n cycles without read signal
    variable read_tb_timeout: integer := 500;
    
  begin

    -- Reset CPU on startup
    reset <= '1';
    run_cycle;
    reset <= '0';

    -- Run clock cycles
    -- Exit loop if read timeout expires
    L: while read_tb_timeout > 0 loop
        run_cycle;
        -- Increment timeout if read signal is not set
        IF rd = '0' THEN
            read_tb_timeout := read_tb_timeout - 1;
        END IF;
    end loop;
    
    -- Print a note & finish simulation now
    assert false report "Simulation finished" severity note;
    wait; -- wait forever (stop simulation)

  end process;

end architecture;
